LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY AUTO_PULSE_MOD IS
GENERIC (PERIOD_W : INTEGER := 6666000);
PORT (	 ENTRADA : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		   CLOCK : IN STD_LOGIC;
	     PULSE_W : OUT INTEGER);
END AUTO_PULSE_MOD;

ARCHITECTURE behavior OF AUTO_PULSE_MOD IS

SIGNAL PULSE_W_I: INTEGER := 0;

BEGIN

	PROCESS (CLOCK)
	
	BEGIN
		IF RISING_EDGE(CLOCK) THEN
			PULSE_W_I <= (PERIOD_W/256) * TO_INTEGER (UNSIGNED(ENTRADA));	
		END IF;
	END PROCESS;
	
	PULSE_W <= PULSE_W_I;

END behavior;