 LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY PWM IS
GENERIC (MAX_PERIODO : INTEGER := 10);--66660000);
PORT (	   	    CLK: IN   STD_LOGIC;
		   MAX_DUTY: IN   INTEGER;
		      SAIDA: OUT  STD_LOGIC);
END PWM;

ARCHITECTURE behavior OF PWM IS
	
	SIGNAL   COUNT : INTEGER   := 0;
	SIGNAL   CLK1  : STD_LOGIC := '0';
	
	BEGIN
	PROCESS (clk)
	BEGIN  
		IF (RISING_EDGE(CLK)) THEN
			COUNT <= COUNT + 1;
			IF (COUNT >= MAX_PERIODO - 1) THEN
				IF (MAX_DUTY <= 0) THEN
					CLK1 <= '0';
				ELSIF (MAX_DUTY >= MAX_PERIODO) THEN
					CLK1 <='1';
				ELSE 
					CLK1 <='1';
				END IF;
				COUNT <= 0;	
			ELSIF (COUNT >= MAX_DUTY - 1) THEN
					CLK1 <= '0';
			END IF;
		END IF;
	END PROCESS;

	
	SAIDA <= CLK1;

END behavior;